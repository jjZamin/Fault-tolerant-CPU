library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity ROMz is
      generic (
                ROM_BYTES : natural := 4000;
                INSTRUCTION_WIDTH : natural := 32;
                DATA_WIDTH : natural := 8;
                ADDR_WIDTH : natural := 32
      );
      Port (
                addr : in std_logic_vector(ADDR_WIDTH - 1 downto 0);
                data_out : out std_logic_vector(INSTRUCTION_WIDTH - 1 downto 0)
      );
end ROMz;

architecture Behavioral of ROMz is
    type ROM_TYPE is array(0 to ROM_BYTES - 1) of std_logic_vector(DATA_WIDTH - 1 downto 0);

    signal ROMz :
    ROM_TYPE :=
                (
-----------------------------------------------------
--SCRUB SEQ
"00110111", "00000000", "00000000", "00000000", --0
"00100011", "00100010", "00010000", "00000000", --4
"00100011", "00100100", "00100000", "00000000", --8
"00100011", "00100110", "00110000", "00000000", --12
"00100011", "00101000", "01000000", "00000000", --16
"00100011", "00101010", "01010000", "00000000", --20
"00100011", "00101100", "01100000", "00000000", --24
"00100011", "00101110", "01110000", "00000000", --28
"00100011", "00100000", "10000000", "00000010", --32
"00100011", "00100010", "10010000", "00000010", --36
"00100011", "00100100", "10100000", "00000010", --40
"00100011", "00100110", "10110000", "00000010", --44
"00100011", "00101000", "11000000", "00000010", --48
"00100011", "00101010", "11010000", "00000010", --52
"00100011", "00101100", "11100000", "00000010", --56
"00100011", "00101110", "11110000", "00000010", --60
"00100011", "00100000", "00000000", "00000101", --64
"00100011", "00100010", "00010000", "00000101", --68
"00100011", "00100100", "00100000", "00000101", --72
"00100011", "00100110", "00110000", "00000101", --76
"00100011", "00101000", "01000000", "00000101", --80
"00100011", "00101010", "01010000", "00000101", --84
"00100011", "00101100", "01100000", "00000101", --88
"00100011", "00101110", "01110000", "00000101", --92
"00100011", "00100000", "10000000", "00000111", --96
"00100011", "00100010", "10010000", "00000111", --100
"00100011", "00100100", "10100000", "00000111", --104
"00100011", "00100110", "10110000", "00000111", --108
"00100011", "00101000", "11000000", "00000111", --112
"00100011", "00101010", "11010000", "00000111", --116
"00100011", "00101100", "11100000", "00000111", --120
"00100011", "00101110", "11110000", "00000111", --124
"11110011", "00010000", "00000000", "01000000", --128
"00100011", "00100000", "00010000", "00000000", --132
"00000000", "00000000", "00000000", "00000000", --136
------------------------------------------------------------
-- LOAD REGISTER AFTER SCRUB OR AT THE BEGINNING OF A PROGRAM.
--
"10000011", "00100000", "01000000", "00000000", --140
"00000011", "00100001", "10000000", "00000000", --144
"10000011", "00100001", "11000000", "00000000", --148
"00000011", "00100010", "00000000", "00000001", --152
"10000011", "00100010", "01000000", "00000001", --156
"00000011", "00100011", "10000000", "00000001", --160
"10000011", "00100011", "11000000", "00000001", --164
"00000011", "00100100", "00000000", "00000010", --168
"10000011", "00100100", "01000000", "00000010", --172
"00000011", "00100101", "10000000", "00000010", --176
"10000011", "00100101", "11000000", "00000010", --180
"00000011", "00100110", "00000000", "00000011", --184
"00000011", "00100111", "01000000", "00000011", --188
"10000011", "00100111", "10000000", "00000011", --192
"00000011", "00101000", "11000000", "00000011", --196
"10000011", "00101000", "00000000", "00000100", --200
"00000011", "00101001", "01000000", "00000100", --204
"10000011", "00101001", "10000000", "00000100", --208
"00000011", "00101010", "11000000", "00000100", --212
"10000011", "00101010", "00000000", "00000101", --216
"00000011", "00101011", "01000000", "00000101", --220
"10000011", "00101011", "10000000", "00000101", --224
"00000011", "00101100", "11000000", "00000101", --228
"10000011", "00101100", "00000000", "00000110", --232
"00000011", "00101101", "01000000", "00000110", --236
"10000011", "00101101", "10000000", "00000110", --240
"00000011", "00101110", "11000000", "00000110", --244
"10000011", "00101110", "00000000", "00000111", --248
"00000011", "00101111", "01000000", "00000111", --252
"10000011", "00101111", "00000000", "00000000", --256
"01100111", "10000000", "00001111", "00000000", --260
-----------------------------------------------------------
--PGORAM!! --264
"00010011", "00000000", "00000000", "00000000",
"10010011", "00000010", "10100000", "00000000",
"00010011", "00000011", "11110000", "00000000",
"10010011", "00000011", "01000000", "01011101",
"00010011", "00000100", "00010000", "00000000",
"00100011", "00100110", "01010000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00100011", "00100110", "01100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"01100111", "00000000", "01000000", "00010110",
"00010011", "00000000", "00000000", "00000000",
"00100011", "10100000", "11100001", "00000001",
"00000011", "00101111", "11000000", "00100000",
"00100011", "00101000", "11100000", "11111111",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00000011", "10101111", "00000001", "00000000",
"01100111", "10000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"10010011", "00000010", "10110000", "00001001",
"00010011", "00000011", "10000000", "01110111",
"10110011", "10000011", "01100010", "01000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"10010011", "00000010", "10100000", "00000000",
"00010011", "00000011", "01000000", "00000001",
"10110011", "10000011", "01100010", "01000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"10010011", "00000010", "10100000", "00000000",
"00010011", "00000011", "00000000", "00000000",
"01100011", "10011000", "01100010", "00000000",
"10010011", "00000011", "10100000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00100011", "00100110", "00000000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00010000", "00000000",
"10010011", "00010011", "01000101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"10010011", "00000100", "01000000", "00000000",
"10110011", "00010011", "10010101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00010000", "00000000",
"10010011", "00000101", "00000000", "00000000",
"01100011", "00001000", "00000000", "00000000",
"10010011", "00000011", "10100000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00000000", "00000010",
"00100011", "00100110", "10100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11010000", "00001101",
"10010011", "00000101", "01010000", "00101011",
"10110011", "01000011", "10110101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"10010011", "00000011", "10100000", "00000000",
"10010011", "01000011", "01010101", "00101011",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"01100011", "01011000", "00000000", "00000000",
"10010011", "00000011", "10100000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00000000", "00000010",
"00100011", "00100110", "10100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11110000", "11111111",
"00100011", "00100110", "10100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"01100011", "01011000", "10100000", "00000000",
"10010011", "00000011", "10100000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00000000", "00000010",
"00100011", "00100110", "10100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11000000", "11111111",
"10010011", "01010011", "00010101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"10010011", "01010011", "00010101", "01000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11110000", "11111111",
"01100011", "01001000", "00000101", "00000000",
"10010011", "00000011", "10100000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00000000", "00000010",
"00100011", "00100110", "10100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11110000", "11111111",
"01100011", "01101000", "10100000", "00000000",
"10010011", "00000011", "10100000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00000000", "00000010",
"00100011", "00100110", "10100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00100011", "00100110", "00000000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11110000", "11111111",
"01100011", "01111000", "00000101", "00000000",
"10010011", "00000011", "10100000", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "00000000", "00000010",
"00100011", "00100110", "10100000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11100000", "11111111",
"10010011", "00000101", "11110000", "11111111",
"10110011", "01110011", "10110101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11110000", "11111111",
"10110011", "01110011", "00000101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "10100000", "00000000",
"10010011", "01100011", "00010101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11110000", "11111111",
"10110011", "01100011", "00000101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "10100000", "00000000",
"10010011", "00100011", "10110101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"00010011", "00000101", "11110000", "11111111",
"10010011", "00000101", "00000000", "00000000",
"10110011", "00110011", "10110101", "00000000",
"00100011", "00100110", "01110000", "00100000",
"11100111", "00000000", "01000000", "00010100",
"00010011", "00000000", "00000000", "00000000",
"01100111", "00000000", "01000000", "00111111",
"00010011", "00000000", "00000000", "00000000",
-----------------------------------------------------------

                    others => x"00"
                );

 attribute rom_style : string;
 attribute rom_style of ROMz : signal is "block";

begin

    data_out(7 downto 0) <= ROMz(to_integer(unsigned(addr)));
    data_out(15 downto 8) <= ROMz(to_integer(unsigned(addr)) + 1);
    data_out(23 downto 16) <= ROMz(to_integer(unsigned(addr)) + 2);
    data_out(31 downto 24) <= ROMz(to_integer(unsigned(addr)) + 3);

end Behavioral;
