library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package SSD1331_ascii_pkg is
  component SSD1331_ascii
        Port (
                  clk : in std_logic;
                  clear : in std_logic;
                  cmd : in std_logic_vector(23 downto 0);
                  addr : in std_logic_vector(31 downto 0);
                  we : in std_logic;
                  SPI_IS_BUSY : in std_logic;

                  spi_addr : out std_logic_vector(31 downto 0);
                  spi_data : out std_logic_vector(7 downto 0);
                  spi_we : out std_logic;
                  ssd_dc : out std_logic;
                  ascii_stall_cpu : out std_logic
        );
  end component;

constant THIS_ADDR : std_logic_vector(31 downto 0) := x"fffffffd";

-- ROM
constant SPI_ADDR_s : std_logic_vector(31 downto 0) := (others => '1');
-- cmds to SSD1331
constant SET_COL_ADDR : std_logic_vector(7 downto 0) := "00010101"; -- x"15";
constant SET_ROW_ADDR : std_logic_vector(7 downto 0) := "01110101"; --x"75";
-- screen size
constant WIDTH : std_logic_vector(7 downto 0) := "01011111";
constant HEIGHT : std_logic_vector(7 downto 0) := "00111111";

-- pix
-- colors [CCCCCBBBBBBAAAAA] -- BGR: first send MSBT, then LSBT
constant WHITE_PIX : std_logic_vector(7 downto 0) := "11111111";
constant BLACK_PIX : std_logic_vector(7 downto 0) := "00000000";

type ROM_TYPE_ascii is array(0 to 3500) of std_logic_vector(7 downto 0); -- 0 to 9
constant ASCII_ROM :
ROM_TYPE_ascii :=
(                            --####################################### 0
                BLACK_PIX, -- 0
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --16
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --32
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --48
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --64
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,--80
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --96
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --112
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, -- 127

                --####################################### 1
                BLACK_PIX, -- 128
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 144
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 160
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 176
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 192
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 208
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 224
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 240
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX, -- 255

                --####################################### 2

                BLACK_PIX, -- 256
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 272
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 288
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 304
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 320
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 336
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 352
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 368
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,  -- 383

                --################################### 3
                BLACK_PIX, -- 384
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 400
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 416
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 432
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 448
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 464
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 480
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 496
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --511

                --################################### 4
                BLACK_PIX, -- 512
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 528
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 544
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 560
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 576
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 592
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 608
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 624
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX, -- 639

                --####################################### 5
                BLACK_PIX, -- 640
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 656
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 672
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 688
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 704
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 720
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 736
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 752
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX, --767

                --##################################### 6

                BLACK_PIX, -- 768
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 784
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 800
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --816
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --832
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --848
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --864
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --880
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,  --895

                --################################## 7

                BLACK_PIX, --896
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --912
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --928
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --944
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,

                BLACK_PIX, --960
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --976
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --992
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1008
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,  --1023

                --################################# 8
                BLACK_PIX, -- 1024
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1040
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1056
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 1072
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1088
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1104
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1120
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1136
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,   -- 1151

                --########################## 9
                BLACK_PIX, -- 1152
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1168
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1184
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1200
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 1216
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1232
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, --1248
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 1264
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                --###################### ALHPABET #######################

                --######################## A

                BLACK_PIX, -- 1264
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                --####################### B
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                --###### C
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                 BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                -- ######## D
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                --####################### E
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                 --####################### F
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                -- ########### R
                BLACK_PIX, -- 1264
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,                

                -- ########### I
                BLACK_PIX, -- 1264
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, 
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,


            --####################################### S
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, 
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 672
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, 
                BLACK_PIX,
                BLACK_PIX, 
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, -- 704
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, 
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, 
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX, 
                BLACK_PIX,
                BLACK_PIX, 
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
              --####################################### V
                BLACK_PIX, -- 0
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX, --16
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX, --32
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX, --48
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX, --64
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX,--80
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX, --96
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX, --96
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                --####################### -
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,

              --####################################### smile
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                
                BLACK_PIX, --96
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,
                
                BLACK_PIX, --96
                BLACK_PIX,
                BLACK_PIX, --96
                BLACK_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                WHITE_PIX,
                BLACK_PIX,
                BLACK_PIX,  
                BLACK_PIX,
                BLACK_PIX,               
                
                 
                others => x"00"
);


 
end package SSD1331_ascii_pkg;
